`timescale 1 ns/10 ps

module bnn_chip(clk,rst,vecY,vecT);
   parameter IWITH = 784;
   parameter OWIDTH = 10;
   parameter NSAMPLES = 10;
   parameter MWIDTH = 4;
   parameter DEPTH = 2;
   input clk,rst
   output reg[OWIDTH:0] vecY, vcT;

   reg[IWIDTH-1:0] vecX;
   reg[MWIDTH-1:0] data_count;

   reg[IWIDTH-1:0] vecXs[0:NSAMPLES-1];
   reg[OWIDTH-1:0] vecTs[0:NSAMPLES-1];

   initial begin
       vecXs[0] = 784'b0000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000001110000000000000000000000000111000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000000100000000000000000000000001110000111000000000000000000110000111110000000000000000111000111111100000000000000011100111101110000000000000001100111000111000000000000001110111000011000000000000000111111100011100000000000000011111100011100000000000000001111111111100000000000000000011111111100000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      vecXs[1] = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000111000011111100000000000000111111111110000000000000000111111100000000000000000000110000000000000000000000000111000000000000000000000000001110000000000000000000000000011110000000000000000000000000011100000000000000000000000000110000000000000000001100000001100000000000000000011111000110000000000000000000111111110000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      vecXs[2] = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000001111000000001000000000000000111000000001100000000000000111000000000110000000000000011100000000011000000000000001100000000001100000000000000111000000001100000000000000111110110000110000000000000001111111110011000000000000000001111111111100000000000000000001101111110000000000000000000000001111000000000000000000000000111100000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000001100000000000000000000000000110000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000;
      vecXs[3] = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000011111111111000000000000000001110000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000001110000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000;
      vecXs[4] = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000111111111111100000000000000011000000001111000000000000000000000000001100000000000000000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000011111100000000000000000001111111000000000000000000011111111000000000000000000000000011000000000000000000000000011100000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000;
      vecXs[5] = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000111111100000000000000000000011111111111000000000000000011111111111110000000000000001111111110111100000000000001111111000001110000000000000111011000000111000000000000011100000000011100000000000011110000000001110000000000001110000000000011000000000000111000000000001100000000000111100000000001110000000000011110000000000111000000000000111000000000011100000000000011110000000011100000000000001111000000011110000000000000011110000011110000000000000001111111111110000000000000000011111111110000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      vecXs[6] = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000111111111111000000000000001111000000001100000000000000110000000000110000000000000011000000000111000000000000001110000000111000000000000000011000000111000000000000000000110000111000000000000000000001100111000000000000000000000111111000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111100000000000000000000001110011000000000000000000000110001100000000000000000000111000111000000000000000000011000011100000000000000000011100000110000000000000000001110000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      vecXs[7] = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111010000000000000000000111111111100000000000000000111100011111000000000000000111100000111000000000000000011000000011110000000000000011100000011110000000000000001100000011110000000000000000110000011110000000000000000011111111110000000000000000001111111110000000000000000000001101110000000000000000000000001110000000000000000000000001111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000;
      vecXs[8] = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000011111111111111110000000000001111111111111110000000000000011111111111100000000000000000111111111000000000000000000001111111110000000000000000001111111111000000000000000000111111111110000000000000000001111001111000000000000000000110000011100000000000000000000000001110000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000011000000111100000000000000011110001111100000000000000001111011111110000000000000000111111111110000000000000000001111111100000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000;
      vecXs[9] = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000111111100000000000000000000111111111100000000000000000001111101111000000000000000000000000011100000000000000000000000001110000000000000000000000000111100000000000000000000000011100000000000000000000000001110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111110000000000000000000000111110000000000000000000000011110000000000000000000000011100000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000;

      vecTs[0] = 10'b0000001000;
      vecTs[1] = 10'b0000010000;
      vecTs[2] = 10'b0000100000;
      vecTs[3] = 10'b0100000000;
      vecTs[4] = 10'b0000100000;
      vecTs[5] = 10'b0000100000;
      vecTs[6] = 10'b0000010000;
      vecTs[7] = 10'b0000100000;
      vecTs[8] = 10'b0001000000;
      vecTs[9] = 10'b0000100000;
   end

   always @(posedge clk) begin
       if (rst == 1) begin
           data_count <= 0;
           vecX <= 0;
           vecT <= 0;
       end
       else begin
           if (data_count < ndata)
               vecX <= vecXs[data_count];
           if (data_count < ndata + DEPTH) begin
               data_count <= data_count + 1;
               vecT <= vectTs[data_count;
           end
           else data_count <= 0;
       end
   end

endmodule
